
entity testbench is

end entity;

architecture TB of testbench is

end architecture;