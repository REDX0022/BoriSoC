arch thing is thing